// audio_nios.v

// Generated using ACDS version 13.1 162 at 2013.12.13.14:52:24

`timescale 1 ps / 1 ps
module audio_nios (
		output wire        c0_out_clk_clk,                             //                  c0_out_clk.clk
		output wire        c0_001_out_clk_clk,                         //              c0_001_out_clk.clk
		input  wire [3:0]  key_external_connection_export,             //     key_external_connection.export
		output wire [3:0]  pio_0_external_connection_export,           //   pio_0_external_connection.export
		input  wire [3:0]  sw_external_connection_export,              //      sw_external_connection.export
		output wire        i2c_scl_external_connection_export,         // i2c_scl_external_connection.export
		inout  wire        i2c_sda_external_connection_export,         // i2c_sda_external_connection.export
		output wire        audio_conduit_end_XCK,                      //           audio_conduit_end.XCK
		input  wire        audio_conduit_end_ADCDAT,                   //                            .ADCDAT
		input  wire        audio_conduit_end_ADCLRC,                   //                            .ADCLRC
		output wire        audio_conduit_end_DACDAT,                   //                            .DACDAT
		input  wire        audio_conduit_end_DACLRC,                   //                            .DACLRC
		input  wire        audio_conduit_end_BCLK,                     //                            .BCLK
		input  wire        clk_clk,                                    //                         clk.clk
		input  wire        reset_reset_n,                              //                       reset.reset_n
		output wire        c2_out_clk_clk,                             //                  c2_out_clk.clk
		output wire [14:0] memory_mem_a,                               //                      memory.mem_a
		output wire [2:0]  memory_mem_ba,                              //                            .mem_ba
		output wire [0:0]  memory_mem_ck,                              //                            .mem_ck
		output wire [0:0]  memory_mem_ck_n,                            //                            .mem_ck_n
		output wire [0:0]  memory_mem_cke,                             //                            .mem_cke
		output wire [0:0]  memory_mem_cs_n,                            //                            .mem_cs_n
		output wire [3:0]  memory_mem_dm,                              //                            .mem_dm
		output wire [0:0]  memory_mem_ras_n,                           //                            .mem_ras_n
		output wire [0:0]  memory_mem_cas_n,                           //                            .mem_cas_n
		output wire [0:0]  memory_mem_we_n,                            //                            .mem_we_n
		output wire        memory_mem_reset_n,                         //                            .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                              //                            .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                             //                            .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                           //                            .mem_dqs_n
		output wire [0:0]  memory_mem_odt,                             //                            .mem_odt
		input  wire        oct_rzqin,                                  //                         oct.rzqin
		output wire        ddr3_status_local_init_done,                //                 ddr3_status.local_init_done
		output wire        ddr3_status_local_cal_success,              //                            .local_cal_success
		output wire        ddr3_status_local_cal_fail,                 //                            .local_cal_fail
		output wire        ddr3_pll_sharing_pll_mem_clk,               //            ddr3_pll_sharing.pll_mem_clk
		output wire        ddr3_pll_sharing_pll_write_clk,             //                            .pll_write_clk
		output wire        ddr3_pll_sharing_pll_locked,                //                            .pll_locked
		output wire        ddr3_pll_sharing_pll_write_clk_pre_phy_clk, //                            .pll_write_clk_pre_phy_clk
		output wire        ddr3_pll_sharing_pll_addr_cmd_clk,          //                            .pll_addr_cmd_clk
		output wire        ddr3_pll_sharing_pll_avl_clk,               //                            .pll_avl_clk
		output wire        ddr3_pll_sharing_pll_config_clk,            //                            .pll_config_clk
		output wire        ddr3_pll_sharing_pll_dr_clk,                //                            .pll_dr_clk
		output wire        ddr3_pll_sharing_pll_dr_clk_pre_phy_clk,    //                            .pll_dr_clk_pre_phy_clk
		output wire        ddr3_pll_sharing_pll_mem_phy_clk,           //                            .pll_mem_phy_clk
		output wire        ddr3_pll_sharing_afi_phy_clk,               //                            .afi_phy_clk
		output wire        ddr3_pll_sharing_pll_avl_phy_clk,           //                            .pll_avl_phy_clk
		input  wire        spi_temperature_external_MISO,              //    spi_temperature_external.MISO
		output wire        spi_temperature_external_MOSI,              //                            .MOSI
		output wire        spi_temperature_external_SCLK,              //                            .SCLK
		output wire        spi_temperature_external_SS_n               //                            .SS_n
	);

	wire          mm_interconnect_0_cpu_peripheral_bridge_s0_waitrequest;        // cpu_peripheral_bridge:s0_waitrequest -> mm_interconnect_0:cpu_peripheral_bridge_s0_waitrequest
	wire    [0:0] mm_interconnect_0_cpu_peripheral_bridge_s0_burstcount;         // mm_interconnect_0:cpu_peripheral_bridge_s0_burstcount -> cpu_peripheral_bridge:s0_burstcount
	wire   [31:0] mm_interconnect_0_cpu_peripheral_bridge_s0_writedata;          // mm_interconnect_0:cpu_peripheral_bridge_s0_writedata -> cpu_peripheral_bridge:s0_writedata
	wire    [8:0] mm_interconnect_0_cpu_peripheral_bridge_s0_address;            // mm_interconnect_0:cpu_peripheral_bridge_s0_address -> cpu_peripheral_bridge:s0_address
	wire          mm_interconnect_0_cpu_peripheral_bridge_s0_write;              // mm_interconnect_0:cpu_peripheral_bridge_s0_write -> cpu_peripheral_bridge:s0_write
	wire          mm_interconnect_0_cpu_peripheral_bridge_s0_read;               // mm_interconnect_0:cpu_peripheral_bridge_s0_read -> cpu_peripheral_bridge:s0_read
	wire   [31:0] mm_interconnect_0_cpu_peripheral_bridge_s0_readdata;           // cpu_peripheral_bridge:s0_readdata -> mm_interconnect_0:cpu_peripheral_bridge_s0_readdata
	wire          mm_interconnect_0_cpu_peripheral_bridge_s0_debugaccess;        // mm_interconnect_0:cpu_peripheral_bridge_s0_debugaccess -> cpu_peripheral_bridge:s0_debugaccess
	wire          mm_interconnect_0_cpu_peripheral_bridge_s0_readdatavalid;      // cpu_peripheral_bridge:s0_readdatavalid -> mm_interconnect_0:cpu_peripheral_bridge_s0_readdatavalid
	wire    [3:0] mm_interconnect_0_cpu_peripheral_bridge_s0_byteenable;         // mm_interconnect_0:cpu_peripheral_bridge_s0_byteenable -> cpu_peripheral_bridge:s0_byteenable
	wire          mm_interconnect_0_cpu_jtag_debug_module_waitrequest;           // cpu:jtag_debug_module_waitrequest -> mm_interconnect_0:cpu_jtag_debug_module_waitrequest
	wire   [31:0] mm_interconnect_0_cpu_jtag_debug_module_writedata;             // mm_interconnect_0:cpu_jtag_debug_module_writedata -> cpu:jtag_debug_module_writedata
	wire    [8:0] mm_interconnect_0_cpu_jtag_debug_module_address;               // mm_interconnect_0:cpu_jtag_debug_module_address -> cpu:jtag_debug_module_address
	wire          mm_interconnect_0_cpu_jtag_debug_module_write;                 // mm_interconnect_0:cpu_jtag_debug_module_write -> cpu:jtag_debug_module_write
	wire          mm_interconnect_0_cpu_jtag_debug_module_read;                  // mm_interconnect_0:cpu_jtag_debug_module_read -> cpu:jtag_debug_module_read
	wire   [31:0] mm_interconnect_0_cpu_jtag_debug_module_readdata;              // cpu:jtag_debug_module_readdata -> mm_interconnect_0:cpu_jtag_debug_module_readdata
	wire          mm_interconnect_0_cpu_jtag_debug_module_debugaccess;           // mm_interconnect_0:cpu_jtag_debug_module_debugaccess -> cpu:jtag_debug_module_debugaccess
	wire    [3:0] mm_interconnect_0_cpu_jtag_debug_module_byteenable;            // mm_interconnect_0:cpu_jtag_debug_module_byteenable -> cpu:jtag_debug_module_byteenable
	wire          mm_interconnect_0_ddr3_avl_waitrequest;                        // DDR3:avl_ready -> mm_interconnect_0:DDR3_avl_waitrequest
	wire    [5:0] mm_interconnect_0_ddr3_avl_burstcount;                         // mm_interconnect_0:DDR3_avl_burstcount -> DDR3:avl_size
	wire  [127:0] mm_interconnect_0_ddr3_avl_writedata;                          // mm_interconnect_0:DDR3_avl_writedata -> DDR3:avl_wdata
	wire   [23:0] mm_interconnect_0_ddr3_avl_address;                            // mm_interconnect_0:DDR3_avl_address -> DDR3:avl_addr
	wire          mm_interconnect_0_ddr3_avl_write;                              // mm_interconnect_0:DDR3_avl_write -> DDR3:avl_write_req
	wire          mm_interconnect_0_ddr3_avl_beginbursttransfer;                 // mm_interconnect_0:DDR3_avl_beginbursttransfer -> DDR3:avl_burstbegin
	wire          mm_interconnect_0_ddr3_avl_read;                               // mm_interconnect_0:DDR3_avl_read -> DDR3:avl_read_req
	wire  [127:0] mm_interconnect_0_ddr3_avl_readdata;                           // DDR3:avl_rdata -> mm_interconnect_0:DDR3_avl_readdata
	wire          mm_interconnect_0_ddr3_avl_readdatavalid;                      // DDR3:avl_rdata_valid -> mm_interconnect_0:DDR3_avl_readdatavalid
	wire   [15:0] mm_interconnect_0_ddr3_avl_byteenable;                         // mm_interconnect_0:DDR3_avl_byteenable -> DDR3:avl_be
	wire   [31:0] mm_interconnect_0_onchip_memory2_1_s1_writedata;               // mm_interconnect_0:onchip_memory2_1_s1_writedata -> onchip_memory2_1:writedata
	wire   [15:0] mm_interconnect_0_onchip_memory2_1_s1_address;                 // mm_interconnect_0:onchip_memory2_1_s1_address -> onchip_memory2_1:address
	wire          mm_interconnect_0_onchip_memory2_1_s1_chipselect;              // mm_interconnect_0:onchip_memory2_1_s1_chipselect -> onchip_memory2_1:chipselect
	wire          mm_interconnect_0_onchip_memory2_1_s1_clken;                   // mm_interconnect_0:onchip_memory2_1_s1_clken -> onchip_memory2_1:clken
	wire          mm_interconnect_0_onchip_memory2_1_s1_write;                   // mm_interconnect_0:onchip_memory2_1_s1_write -> onchip_memory2_1:write
	wire   [31:0] mm_interconnect_0_onchip_memory2_1_s1_readdata;                // onchip_memory2_1:readdata -> mm_interconnect_0:onchip_memory2_1_s1_readdata
	wire    [3:0] mm_interconnect_0_onchip_memory2_1_s1_byteenable;              // mm_interconnect_0:onchip_memory2_1_s1_byteenable -> onchip_memory2_1:byteenable
	wire          cpu_instruction_master_waitrequest;                            // mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	wire   [28:0] cpu_instruction_master_address;                                // cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	wire          cpu_instruction_master_read;                                   // cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	wire   [31:0] cpu_instruction_master_readdata;                               // mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	wire          cpu_instruction_master_readdatavalid;                          // mm_interconnect_0:cpu_instruction_master_readdatavalid -> cpu:i_readdatavalid
	wire   [15:0] mm_interconnect_0_audio_avalon_slave_writedata;                // mm_interconnect_0:audio_avalon_slave_writedata -> audio:avs_s1_writedata
	wire    [2:0] mm_interconnect_0_audio_avalon_slave_address;                  // mm_interconnect_0:audio_avalon_slave_address -> audio:avs_s1_address
	wire          mm_interconnect_0_audio_avalon_slave_write;                    // mm_interconnect_0:audio_avalon_slave_write -> audio:avs_s1_write
	wire          mm_interconnect_0_audio_avalon_slave_read;                     // mm_interconnect_0:audio_avalon_slave_read -> audio:avs_s1_read
	wire   [15:0] mm_interconnect_0_audio_avalon_slave_readdata;                 // audio:avs_s1_readdata -> mm_interconnect_0:audio_avalon_slave_readdata
	wire          mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest;     // jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	wire   [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata;       // mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	wire    [0:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_address;         // mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	wire          mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect;      // mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	wire          mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;           // mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> jtag_uart:av_write_n
	wire          mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;            // mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> jtag_uart:av_read_n
	wire   [31:0] mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata;        // jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	wire          ddr3_afi_clk_clk;                                              // DDR3:afi_clk -> [mm_interconnect_0:DDR3_afi_clk_clk, rst_controller_009:clk]
	wire   [15:0] mm_interconnect_0_timer_s1_writedata;                          // mm_interconnect_0:timer_s1_writedata -> timer:writedata
	wire    [2:0] mm_interconnect_0_timer_s1_address;                            // mm_interconnect_0:timer_s1_address -> timer:address
	wire          mm_interconnect_0_timer_s1_chipselect;                         // mm_interconnect_0:timer_s1_chipselect -> timer:chipselect
	wire          mm_interconnect_0_timer_s1_write;                              // mm_interconnect_0:timer_s1_write -> timer:write_n
	wire   [15:0] mm_interconnect_0_timer_s1_readdata;                           // timer:readdata -> mm_interconnect_0:timer_s1_readdata
	wire          cpu_data_master_waitrequest;                                   // mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	wire   [31:0] cpu_data_master_writedata;                                     // cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	wire   [28:0] cpu_data_master_address;                                       // cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	wire          cpu_data_master_write;                                         // cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	wire          cpu_data_master_read;                                          // cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	wire   [31:0] cpu_data_master_readdata;                                      // mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	wire          cpu_data_master_debugaccess;                                   // cpu:jtag_debug_module_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	wire          cpu_data_master_readdatavalid;                                 // mm_interconnect_0:cpu_data_master_readdatavalid -> cpu:d_readdatavalid
	wire    [3:0] cpu_data_master_byteenable;                                    // cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	wire   [15:0] mm_interconnect_0_spi_temperature_spi_control_port_writedata;  // mm_interconnect_0:spi_temperature_spi_control_port_writedata -> spi_temperature:data_from_cpu
	wire    [2:0] mm_interconnect_0_spi_temperature_spi_control_port_address;    // mm_interconnect_0:spi_temperature_spi_control_port_address -> spi_temperature:mem_addr
	wire          mm_interconnect_0_spi_temperature_spi_control_port_chipselect; // mm_interconnect_0:spi_temperature_spi_control_port_chipselect -> spi_temperature:spi_select
	wire          mm_interconnect_0_spi_temperature_spi_control_port_write;      // mm_interconnect_0:spi_temperature_spi_control_port_write -> spi_temperature:write_n
	wire          mm_interconnect_0_spi_temperature_spi_control_port_read;       // mm_interconnect_0:spi_temperature_spi_control_port_read -> spi_temperature:read_n
	wire   [15:0] mm_interconnect_0_spi_temperature_spi_control_port_readdata;   // spi_temperature:data_to_cpu -> mm_interconnect_0:spi_temperature_spi_control_port_readdata
	wire    [0:0] mm_interconnect_0_sysid_qsys_control_slave_address;            // mm_interconnect_0:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire   [31:0] mm_interconnect_0_sysid_qsys_control_slave_readdata;           // sysid_qsys:readdata -> mm_interconnect_0:sysid_qsys_control_slave_readdata
	wire   [31:0] mm_interconnect_1_sw_s1_writedata;                             // mm_interconnect_1:sw_s1_writedata -> sw:writedata
	wire    [1:0] mm_interconnect_1_sw_s1_address;                               // mm_interconnect_1:sw_s1_address -> sw:address
	wire          mm_interconnect_1_sw_s1_chipselect;                            // mm_interconnect_1:sw_s1_chipselect -> sw:chipselect
	wire          mm_interconnect_1_sw_s1_write;                                 // mm_interconnect_1:sw_s1_write -> sw:write_n
	wire   [31:0] mm_interconnect_1_sw_s1_readdata;                              // sw:readdata -> mm_interconnect_1:sw_s1_readdata
	wire   [31:0] mm_interconnect_1_key_s1_writedata;                            // mm_interconnect_1:key_s1_writedata -> key:writedata
	wire    [1:0] mm_interconnect_1_key_s1_address;                              // mm_interconnect_1:key_s1_address -> key:address
	wire          mm_interconnect_1_key_s1_chipselect;                           // mm_interconnect_1:key_s1_chipselect -> key:chipselect
	wire          mm_interconnect_1_key_s1_write;                                // mm_interconnect_1:key_s1_write -> key:write_n
	wire   [31:0] mm_interconnect_1_key_s1_readdata;                             // key:readdata -> mm_interconnect_1:key_s1_readdata
	wire   [31:0] mm_interconnect_1_i2c_scl_s1_writedata;                        // mm_interconnect_1:i2c_scl_s1_writedata -> i2c_scl:writedata
	wire    [1:0] mm_interconnect_1_i2c_scl_s1_address;                          // mm_interconnect_1:i2c_scl_s1_address -> i2c_scl:address
	wire          mm_interconnect_1_i2c_scl_s1_chipselect;                       // mm_interconnect_1:i2c_scl_s1_chipselect -> i2c_scl:chipselect
	wire          mm_interconnect_1_i2c_scl_s1_write;                            // mm_interconnect_1:i2c_scl_s1_write -> i2c_scl:write_n
	wire   [31:0] mm_interconnect_1_i2c_scl_s1_readdata;                         // i2c_scl:readdata -> mm_interconnect_1:i2c_scl_s1_readdata
	wire    [0:0] cpu_peripheral_bridge_m0_burstcount;                           // cpu_peripheral_bridge:m0_burstcount -> mm_interconnect_1:cpu_peripheral_bridge_m0_burstcount
	wire          cpu_peripheral_bridge_m0_waitrequest;                          // mm_interconnect_1:cpu_peripheral_bridge_m0_waitrequest -> cpu_peripheral_bridge:m0_waitrequest
	wire    [8:0] cpu_peripheral_bridge_m0_address;                              // cpu_peripheral_bridge:m0_address -> mm_interconnect_1:cpu_peripheral_bridge_m0_address
	wire   [31:0] cpu_peripheral_bridge_m0_writedata;                            // cpu_peripheral_bridge:m0_writedata -> mm_interconnect_1:cpu_peripheral_bridge_m0_writedata
	wire          cpu_peripheral_bridge_m0_write;                                // cpu_peripheral_bridge:m0_write -> mm_interconnect_1:cpu_peripheral_bridge_m0_write
	wire          cpu_peripheral_bridge_m0_read;                                 // cpu_peripheral_bridge:m0_read -> mm_interconnect_1:cpu_peripheral_bridge_m0_read
	wire   [31:0] cpu_peripheral_bridge_m0_readdata;                             // mm_interconnect_1:cpu_peripheral_bridge_m0_readdata -> cpu_peripheral_bridge:m0_readdata
	wire          cpu_peripheral_bridge_m0_debugaccess;                          // cpu_peripheral_bridge:m0_debugaccess -> mm_interconnect_1:cpu_peripheral_bridge_m0_debugaccess
	wire    [3:0] cpu_peripheral_bridge_m0_byteenable;                           // cpu_peripheral_bridge:m0_byteenable -> mm_interconnect_1:cpu_peripheral_bridge_m0_byteenable
	wire          cpu_peripheral_bridge_m0_readdatavalid;                        // mm_interconnect_1:cpu_peripheral_bridge_m0_readdatavalid -> cpu_peripheral_bridge:m0_readdatavalid
	wire   [31:0] mm_interconnect_1_pio_led_s1_writedata;                        // mm_interconnect_1:pio_led_s1_writedata -> pio_led:writedata
	wire    [1:0] mm_interconnect_1_pio_led_s1_address;                          // mm_interconnect_1:pio_led_s1_address -> pio_led:address
	wire          mm_interconnect_1_pio_led_s1_chipselect;                       // mm_interconnect_1:pio_led_s1_chipselect -> pio_led:chipselect
	wire          mm_interconnect_1_pio_led_s1_write;                            // mm_interconnect_1:pio_led_s1_write -> pio_led:write_n
	wire   [31:0] mm_interconnect_1_pio_led_s1_readdata;                         // pio_led:readdata -> mm_interconnect_1:pio_led_s1_readdata
	wire   [31:0] mm_interconnect_1_i2c_sda_s1_writedata;                        // mm_interconnect_1:i2c_sda_s1_writedata -> i2c_sda:writedata
	wire    [1:0] mm_interconnect_1_i2c_sda_s1_address;                          // mm_interconnect_1:i2c_sda_s1_address -> i2c_sda:address
	wire          mm_interconnect_1_i2c_sda_s1_chipselect;                       // mm_interconnect_1:i2c_sda_s1_chipselect -> i2c_sda:chipselect
	wire          mm_interconnect_1_i2c_sda_s1_write;                            // mm_interconnect_1:i2c_sda_s1_write -> i2c_sda:write_n
	wire   [31:0] mm_interconnect_1_i2c_sda_s1_readdata;                         // i2c_sda:readdata -> mm_interconnect_1:i2c_sda_s1_readdata
	wire          irq_mapper_receiver0_irq;                                      // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire   [31:0] cpu_d_irq_irq;                                                 // irq_mapper:sender_irq -> cpu:d_irq
	wire          irq_mapper_receiver1_irq;                                      // irq_synchronizer:sender_irq -> irq_mapper:receiver1_irq
	wire    [0:0] irq_synchronizer_receiver_irq;                                 // key:irq -> irq_synchronizer:receiver_irq
	wire          irq_mapper_receiver2_irq;                                      // irq_synchronizer_001:sender_irq -> irq_mapper:receiver2_irq
	wire    [0:0] irq_synchronizer_001_receiver_irq;                             // sw:irq -> irq_synchronizer_001:receiver_irq
	wire          irq_mapper_receiver3_irq;                                      // irq_synchronizer_002:sender_irq -> irq_mapper:receiver3_irq
	wire    [0:0] irq_synchronizer_002_receiver_irq;                             // timer:irq -> irq_synchronizer_002:receiver_irq
	wire          irq_mapper_receiver4_irq;                                      // irq_synchronizer_003:sender_irq -> irq_mapper:receiver4_irq
	wire    [0:0] irq_synchronizer_003_receiver_irq;                             // spi_temperature:irq -> irq_synchronizer_003:receiver_irq
	wire          rst_controller_reset_out_reset;                                // rst_controller:reset_out -> [cpu_peripheral_bridge:m0_reset, mm_interconnect_1:cpu_peripheral_bridge_m0_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_001_reset_out_reset;                            // rst_controller_001:reset_out -> [cpu_peripheral_bridge:s0_reset, mm_interconnect_0:cpu_peripheral_bridge_s0_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_002_reset_out_reset;                            // rst_controller_002:reset_out -> [cpu:reset_n, irq_mapper:reset, irq_synchronizer:sender_reset, irq_synchronizer_001:sender_reset, irq_synchronizer_002:sender_reset, irq_synchronizer_003:sender_reset, jtag_uart:rst_n, mm_interconnect_0:cpu_reset_n_reset_bridge_in_reset_reset, onchip_memory2_1:reset, rst_translator:in_reset]
	wire          rst_controller_002_reset_out_reset_req;                        // rst_controller_002:reset_req -> [cpu:reset_req, onchip_memory2_1:reset_req, rst_translator:reset_req_in]
	wire          cpu_jtag_debug_module_reset_reset;                             // cpu:jtag_debug_module_resetrequest -> [rst_controller_002:reset_in0, rst_controller_003:reset_in0, rst_controller_004:reset_in0, rst_controller_006:reset_in1, rst_controller_007:reset_in1, rst_controller_008:reset_in1]
	wire          rst_controller_003_reset_out_reset;                            // rst_controller_003:reset_out -> [i2c_scl:reset_n, i2c_sda:reset_n, irq_synchronizer:receiver_reset, irq_synchronizer_001:receiver_reset, key:reset_n, mm_interconnect_1:key_reset_reset_bridge_in_reset_reset, pio_led:reset_n, sw:reset_n]
	wire          rst_controller_004_reset_out_reset;                            // rst_controller_004:reset_out -> [audio:avs_s1_reset, mm_interconnect_0:audio_clock_sink_reset_reset_bridge_in_reset_reset]
	wire          rst_controller_005_reset_out_reset;                            // rst_controller_005:reset_out -> [altpll:rst, altpll_audio:rst]
	wire          rst_controller_006_reset_out_reset;                            // rst_controller_006:reset_out -> DDR3:global_reset_n
	wire          rst_controller_007_reset_out_reset;                            // rst_controller_007:reset_out -> DDR3:soft_reset_n
	wire          rst_controller_008_reset_out_reset;                            // rst_controller_008:reset_out -> [irq_synchronizer_002:receiver_reset, irq_synchronizer_003:receiver_reset, mm_interconnect_0:timer_reset_reset_bridge_in_reset_reset, spi_temperature:reset_n, sysid_qsys:reset_n, timer:reset_n]
	wire          rst_controller_009_reset_out_reset;                            // rst_controller_009:reset_out -> mm_interconnect_0:DDR3_avl_translator_reset_reset_bridge_in_reset_reset
	wire          ddr3_afi_reset_reset;                                          // DDR3:afi_reset_n -> rst_controller_009:reset_in0

	altera_avalon_mm_clock_crossing_bridge #(
		.DATA_WIDTH          (32),
		.SYMBOL_WIDTH        (8),
		.ADDRESS_WIDTH       (9),
		.BURSTCOUNT_WIDTH    (1),
		.COMMAND_FIFO_DEPTH  (32),
		.RESPONSE_FIFO_DEPTH (64),
		.MASTER_SYNC_DEPTH   (3),
		.SLAVE_SYNC_DEPTH    (3)
	) cpu_peripheral_bridge (
		.m0_clk           (c2_out_clk_clk),                                           //   m0_clk.clk
		.m0_reset         (rst_controller_reset_out_reset),                           // m0_reset.reset
		.s0_clk           (c0_001_out_clk_clk),                                       //   s0_clk.clk
		.s0_reset         (rst_controller_001_reset_out_reset),                       // s0_reset.reset
		.s0_waitrequest   (mm_interconnect_0_cpu_peripheral_bridge_s0_waitrequest),   //       s0.waitrequest
		.s0_readdata      (mm_interconnect_0_cpu_peripheral_bridge_s0_readdata),      //         .readdata
		.s0_readdatavalid (mm_interconnect_0_cpu_peripheral_bridge_s0_readdatavalid), //         .readdatavalid
		.s0_burstcount    (mm_interconnect_0_cpu_peripheral_bridge_s0_burstcount),    //         .burstcount
		.s0_writedata     (mm_interconnect_0_cpu_peripheral_bridge_s0_writedata),     //         .writedata
		.s0_address       (mm_interconnect_0_cpu_peripheral_bridge_s0_address),       //         .address
		.s0_write         (mm_interconnect_0_cpu_peripheral_bridge_s0_write),         //         .write
		.s0_read          (mm_interconnect_0_cpu_peripheral_bridge_s0_read),          //         .read
		.s0_byteenable    (mm_interconnect_0_cpu_peripheral_bridge_s0_byteenable),    //         .byteenable
		.s0_debugaccess   (mm_interconnect_0_cpu_peripheral_bridge_s0_debugaccess),   //         .debugaccess
		.m0_waitrequest   (cpu_peripheral_bridge_m0_waitrequest),                     //       m0.waitrequest
		.m0_readdata      (cpu_peripheral_bridge_m0_readdata),                        //         .readdata
		.m0_readdatavalid (cpu_peripheral_bridge_m0_readdatavalid),                   //         .readdatavalid
		.m0_burstcount    (cpu_peripheral_bridge_m0_burstcount),                      //         .burstcount
		.m0_writedata     (cpu_peripheral_bridge_m0_writedata),                       //         .writedata
		.m0_address       (cpu_peripheral_bridge_m0_address),                         //         .address
		.m0_write         (cpu_peripheral_bridge_m0_write),                           //         .write
		.m0_read          (cpu_peripheral_bridge_m0_read),                            //         .read
		.m0_byteenable    (cpu_peripheral_bridge_m0_byteenable),                      //         .byteenable
		.m0_debugaccess   (cpu_peripheral_bridge_m0_debugaccess)                      //         .debugaccess
	);

	audio_nios_cpu cpu (
		.clk                                   (c0_001_out_clk_clk),                                  //                       clk.clk
		.reset_n                               (~rst_controller_002_reset_out_reset),                 //                   reset_n.reset_n
		.reset_req                             (rst_controller_002_reset_out_reset_req),              //                          .reset_req
		.d_address                             (cpu_data_master_address),                             //               data_master.address
		.d_byteenable                          (cpu_data_master_byteenable),                          //                          .byteenable
		.d_read                                (cpu_data_master_read),                                //                          .read
		.d_readdata                            (cpu_data_master_readdata),                            //                          .readdata
		.d_waitrequest                         (cpu_data_master_waitrequest),                         //                          .waitrequest
		.d_write                               (cpu_data_master_write),                               //                          .write
		.d_writedata                           (cpu_data_master_writedata),                           //                          .writedata
		.d_readdatavalid                       (cpu_data_master_readdatavalid),                       //                          .readdatavalid
		.jtag_debug_module_debugaccess_to_roms (cpu_data_master_debugaccess),                         //                          .debugaccess
		.i_address                             (cpu_instruction_master_address),                      //        instruction_master.address
		.i_read                                (cpu_instruction_master_read),                         //                          .read
		.i_readdata                            (cpu_instruction_master_readdata),                     //                          .readdata
		.i_waitrequest                         (cpu_instruction_master_waitrequest),                  //                          .waitrequest
		.i_readdatavalid                       (cpu_instruction_master_readdatavalid),                //                          .readdatavalid
		.d_irq                                 (cpu_d_irq_irq),                                       //                     d_irq.irq
		.jtag_debug_module_resetrequest        (cpu_jtag_debug_module_reset_reset),                   //   jtag_debug_module_reset.reset
		.jtag_debug_module_address             (mm_interconnect_0_cpu_jtag_debug_module_address),     //         jtag_debug_module.address
		.jtag_debug_module_byteenable          (mm_interconnect_0_cpu_jtag_debug_module_byteenable),  //                          .byteenable
		.jtag_debug_module_debugaccess         (mm_interconnect_0_cpu_jtag_debug_module_debugaccess), //                          .debugaccess
		.jtag_debug_module_read                (mm_interconnect_0_cpu_jtag_debug_module_read),        //                          .read
		.jtag_debug_module_readdata            (mm_interconnect_0_cpu_jtag_debug_module_readdata),    //                          .readdata
		.jtag_debug_module_waitrequest         (mm_interconnect_0_cpu_jtag_debug_module_waitrequest), //                          .waitrequest
		.jtag_debug_module_write               (mm_interconnect_0_cpu_jtag_debug_module_write),       //                          .write
		.jtag_debug_module_writedata           (mm_interconnect_0_cpu_jtag_debug_module_writedata),   //                          .writedata
		.no_ci_readra                          ()                                                     // custom_instruction_master.readra
	);

	audio_nios_jtag_uart jtag_uart (
		.clk            (c0_001_out_clk_clk),                                        //               clk.clk
		.rst_n          (~rst_controller_002_reset_out_reset),                       //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                   //               irq.irq
	);

	audio_nios_key key (
		.clk        (c2_out_clk_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_003_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_1_key_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_key_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_key_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_key_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_key_s1_readdata),   //                    .readdata
		.in_port    (key_external_connection_export),      // external_connection.export
		.irq        (irq_synchronizer_receiver_irq)        //                 irq.irq
	);

	audio_nios_pio_led pio_led (
		.clk        (c2_out_clk_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_003_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_1_pio_led_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_pio_led_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_pio_led_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_pio_led_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_pio_led_s1_readdata),   //                    .readdata
		.out_port   (pio_0_external_connection_export)         // external_connection.export
	);

	audio_nios_key sw (
		.clk        (c2_out_clk_clk),                      //                 clk.clk
		.reset_n    (~rst_controller_003_reset_out_reset), //               reset.reset_n
		.address    (mm_interconnect_1_sw_s1_address),     //                  s1.address
		.write_n    (~mm_interconnect_1_sw_s1_write),      //                    .write_n
		.writedata  (mm_interconnect_1_sw_s1_writedata),   //                    .writedata
		.chipselect (mm_interconnect_1_sw_s1_chipselect),  //                    .chipselect
		.readdata   (mm_interconnect_1_sw_s1_readdata),    //                    .readdata
		.in_port    (sw_external_connection_export),       // external_connection.export
		.irq        (irq_synchronizer_001_receiver_irq)    //                 irq.irq
	);

	audio_nios_i2c_scl i2c_scl (
		.clk        (c2_out_clk_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_003_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_1_i2c_scl_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_i2c_scl_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_i2c_scl_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_i2c_scl_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_i2c_scl_s1_readdata),   //                    .readdata
		.out_port   (i2c_scl_external_connection_export)       // external_connection.export
	);

	audio_nios_i2c_sda i2c_sda (
		.clk        (c2_out_clk_clk),                          //                 clk.clk
		.reset_n    (~rst_controller_003_reset_out_reset),     //               reset.reset_n
		.address    (mm_interconnect_1_i2c_sda_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_1_i2c_sda_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_1_i2c_sda_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_1_i2c_sda_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_1_i2c_sda_s1_readdata),   //                    .readdata
		.bidir_port (i2c_sda_external_connection_export)       // external_connection.export
	);

	audio_nios_audio audio (
		.avs_s1_address       (mm_interconnect_0_audio_avalon_slave_address),   //     avalon_slave.address
		.avs_s1_read          (mm_interconnect_0_audio_avalon_slave_read),      //                 .read
		.avs_s1_readdata      (mm_interconnect_0_audio_avalon_slave_readdata),  //                 .readdata
		.avs_s1_write         (mm_interconnect_0_audio_avalon_slave_write),     //                 .write
		.avs_s1_writedata     (mm_interconnect_0_audio_avalon_slave_writedata), //                 .writedata
		.avs_s1_clk           (c0_out_clk_clk),                                 //       clock_sink.clk
		.avs_s1_reset         (rst_controller_004_reset_out_reset),             // clock_sink_reset.reset
		.avs_s1_export_XCK    (audio_conduit_end_XCK),                          //      conduit_end.export
		.avs_s1_export_ADCDAT (audio_conduit_end_ADCDAT),                       //                 .export
		.avs_s1_export_ADCLRC (audio_conduit_end_ADCLRC),                       //                 .export
		.avs_s1_export_DACDAT (audio_conduit_end_DACDAT),                       //                 .export
		.avs_s1_export_DACLRC (audio_conduit_end_DACLRC),                       //                 .export
		.avs_s1_export_BCLK   (audio_conduit_end_BCLK)                          //                 .export
	);

	audio_nios_onchip_memory2_1 onchip_memory2_1 (
		.clk        (c0_001_out_clk_clk),                               //   clk1.clk
		.address    (mm_interconnect_0_onchip_memory2_1_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_onchip_memory2_1_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_onchip_memory2_1_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_onchip_memory2_1_s1_write),      //       .write
		.readdata   (mm_interconnect_0_onchip_memory2_1_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_onchip_memory2_1_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_onchip_memory2_1_s1_byteenable), //       .byteenable
		.reset      (rst_controller_002_reset_out_reset),               // reset1.reset
		.reset_req  (rst_controller_002_reset_out_reset_req)            //       .reset_req
	);

	audio_nios_altpll_audio altpll_audio (
		.refclk   (clk_clk),                            //  refclk.clk
		.rst      (rst_controller_005_reset_out_reset), //   reset.reset
		.outclk_0 (c0_out_clk_clk),                     // outclk0.clk
		.locked   ()                                    // (terminated)
	);

	audio_nios_altpll altpll (
		.refclk   (clk_clk),                            //  refclk.clk
		.rst      (rst_controller_005_reset_out_reset), //   reset.reset
		.outclk_0 (c0_001_out_clk_clk),                 // outclk0.clk
		.outclk_1 (c2_out_clk_clk),                     // outclk1.clk
		.outclk_2 (),                                   // outclk2.clk
		.locked   ()                                    // (terminated)
	);

	audio_nios_DDR3 ddr3 (
		.pll_ref_clk               (clk_clk),                                       //      pll_ref_clk.clk
		.global_reset_n            (~rst_controller_006_reset_out_reset),           //     global_reset.reset_n
		.soft_reset_n              (~rst_controller_007_reset_out_reset),           //       soft_reset.reset_n
		.afi_clk                   (ddr3_afi_clk_clk),                              //          afi_clk.clk
		.afi_half_clk              (),                                              //     afi_half_clk.clk
		.afi_reset_n               (ddr3_afi_reset_reset),                          //        afi_reset.reset_n
		.afi_reset_export_n        (),                                              // afi_reset_export.reset_n
		.mem_a                     (memory_mem_a),                                  //           memory.mem_a
		.mem_ba                    (memory_mem_ba),                                 //                 .mem_ba
		.mem_ck                    (memory_mem_ck),                                 //                 .mem_ck
		.mem_ck_n                  (memory_mem_ck_n),                               //                 .mem_ck_n
		.mem_cke                   (memory_mem_cke),                                //                 .mem_cke
		.mem_cs_n                  (memory_mem_cs_n),                               //                 .mem_cs_n
		.mem_dm                    (memory_mem_dm),                                 //                 .mem_dm
		.mem_ras_n                 (memory_mem_ras_n),                              //                 .mem_ras_n
		.mem_cas_n                 (memory_mem_cas_n),                              //                 .mem_cas_n
		.mem_we_n                  (memory_mem_we_n),                               //                 .mem_we_n
		.mem_reset_n               (memory_mem_reset_n),                            //                 .mem_reset_n
		.mem_dq                    (memory_mem_dq),                                 //                 .mem_dq
		.mem_dqs                   (memory_mem_dqs),                                //                 .mem_dqs
		.mem_dqs_n                 (memory_mem_dqs_n),                              //                 .mem_dqs_n
		.mem_odt                   (memory_mem_odt),                                //                 .mem_odt
		.avl_ready                 (mm_interconnect_0_ddr3_avl_waitrequest),        //              avl.waitrequest_n
		.avl_burstbegin            (mm_interconnect_0_ddr3_avl_beginbursttransfer), //                 .beginbursttransfer
		.avl_addr                  (mm_interconnect_0_ddr3_avl_address),            //                 .address
		.avl_rdata_valid           (mm_interconnect_0_ddr3_avl_readdatavalid),      //                 .readdatavalid
		.avl_rdata                 (mm_interconnect_0_ddr3_avl_readdata),           //                 .readdata
		.avl_wdata                 (mm_interconnect_0_ddr3_avl_writedata),          //                 .writedata
		.avl_be                    (mm_interconnect_0_ddr3_avl_byteenable),         //                 .byteenable
		.avl_read_req              (mm_interconnect_0_ddr3_avl_read),               //                 .read
		.avl_write_req             (mm_interconnect_0_ddr3_avl_write),              //                 .write
		.avl_size                  (mm_interconnect_0_ddr3_avl_burstcount),         //                 .burstcount
		.local_init_done           (ddr3_status_local_init_done),                   //           status.local_init_done
		.local_cal_success         (ddr3_status_local_cal_success),                 //                 .local_cal_success
		.local_cal_fail            (ddr3_status_local_cal_fail),                    //                 .local_cal_fail
		.oct_rzqin                 (oct_rzqin),                                     //              oct.rzqin
		.pll_mem_clk               (ddr3_pll_sharing_pll_mem_clk),                  //      pll_sharing.pll_mem_clk
		.pll_write_clk             (ddr3_pll_sharing_pll_write_clk),                //                 .pll_write_clk
		.pll_locked                (ddr3_pll_sharing_pll_locked),                   //                 .pll_locked
		.pll_write_clk_pre_phy_clk (ddr3_pll_sharing_pll_write_clk_pre_phy_clk),    //                 .pll_write_clk_pre_phy_clk
		.pll_addr_cmd_clk          (ddr3_pll_sharing_pll_addr_cmd_clk),             //                 .pll_addr_cmd_clk
		.pll_avl_clk               (ddr3_pll_sharing_pll_avl_clk),                  //                 .pll_avl_clk
		.pll_config_clk            (ddr3_pll_sharing_pll_config_clk),               //                 .pll_config_clk
		.pll_dr_clk                (ddr3_pll_sharing_pll_dr_clk),                   //                 .pll_dr_clk
		.pll_dr_clk_pre_phy_clk    (ddr3_pll_sharing_pll_dr_clk_pre_phy_clk),       //                 .pll_dr_clk_pre_phy_clk
		.pll_mem_phy_clk           (ddr3_pll_sharing_pll_mem_phy_clk),              //                 .pll_mem_phy_clk
		.afi_phy_clk               (ddr3_pll_sharing_afi_phy_clk),                  //                 .afi_phy_clk
		.pll_avl_phy_clk           (ddr3_pll_sharing_pll_avl_phy_clk)               //                 .pll_avl_phy_clk
	);

	audio_nios_timer timer (
		.clk        (clk_clk),                               //   clk.clk
		.reset_n    (~rst_controller_008_reset_out_reset),   // reset.reset_n
		.address    (mm_interconnect_0_timer_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timer_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timer_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timer_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timer_s1_write),     //      .write_n
		.irq        (irq_synchronizer_002_receiver_irq)      //   irq.irq
	);

	audio_nios_sysid_qsys sysid_qsys (
		.clock    (clk_clk),                                             //           clk.clk
		.reset_n  (~rst_controller_008_reset_out_reset),                 //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_control_slave_address)   //              .address
	);

	audio_nios_spi_temperature spi_temperature (
		.clk           (clk_clk),                                                       //              clk.clk
		.reset_n       (~rst_controller_008_reset_out_reset),                           //            reset.reset_n
		.data_from_cpu (mm_interconnect_0_spi_temperature_spi_control_port_writedata),  // spi_control_port.writedata
		.data_to_cpu   (mm_interconnect_0_spi_temperature_spi_control_port_readdata),   //                 .readdata
		.mem_addr      (mm_interconnect_0_spi_temperature_spi_control_port_address),    //                 .address
		.read_n        (~mm_interconnect_0_spi_temperature_spi_control_port_read),      //                 .read_n
		.spi_select    (mm_interconnect_0_spi_temperature_spi_control_port_chipselect), //                 .chipselect
		.write_n       (~mm_interconnect_0_spi_temperature_spi_control_port_write),     //                 .write_n
		.irq           (irq_synchronizer_003_receiver_irq),                             //              irq.irq
		.MISO          (spi_temperature_external_MISO),                                 //         external.export
		.MOSI          (spi_temperature_external_MOSI),                                 //                 .export
		.SCLK          (spi_temperature_external_SCLK),                                 //                 .export
		.SS_n          (spi_temperature_external_SS_n)                                  //                 .export
	);

	audio_nios_mm_interconnect_0 mm_interconnect_0 (
		.altpll_outclk0_clk                                         (c0_001_out_clk_clk),                                            //                                       altpll_outclk0.clk
		.altpll_audio_outclk0_clk                                   (c0_out_clk_clk),                                                //                                 altpll_audio_outclk0.clk
		.clk_50_clk_clk                                             (clk_clk),                                                       //                                           clk_50_clk.clk
		.DDR3_afi_clk_clk                                           (ddr3_afi_clk_clk),                                              //                                         DDR3_afi_clk.clk
		.audio_clock_sink_reset_reset_bridge_in_reset_reset         (rst_controller_004_reset_out_reset),                            //         audio_clock_sink_reset_reset_bridge_in_reset.reset
		.cpu_peripheral_bridge_s0_reset_reset_bridge_in_reset_reset (rst_controller_001_reset_out_reset),                            // cpu_peripheral_bridge_s0_reset_reset_bridge_in_reset.reset
		.cpu_reset_n_reset_bridge_in_reset_reset                    (rst_controller_002_reset_out_reset),                            //                    cpu_reset_n_reset_bridge_in_reset.reset
		.DDR3_avl_translator_reset_reset_bridge_in_reset_reset      (rst_controller_009_reset_out_reset),                            //      DDR3_avl_translator_reset_reset_bridge_in_reset.reset
		.timer_reset_reset_bridge_in_reset_reset                    (rst_controller_008_reset_out_reset),                            //                    timer_reset_reset_bridge_in_reset.reset
		.cpu_data_master_address                                    (cpu_data_master_address),                                       //                                      cpu_data_master.address
		.cpu_data_master_waitrequest                                (cpu_data_master_waitrequest),                                   //                                                     .waitrequest
		.cpu_data_master_byteenable                                 (cpu_data_master_byteenable),                                    //                                                     .byteenable
		.cpu_data_master_read                                       (cpu_data_master_read),                                          //                                                     .read
		.cpu_data_master_readdata                                   (cpu_data_master_readdata),                                      //                                                     .readdata
		.cpu_data_master_readdatavalid                              (cpu_data_master_readdatavalid),                                 //                                                     .readdatavalid
		.cpu_data_master_write                                      (cpu_data_master_write),                                         //                                                     .write
		.cpu_data_master_writedata                                  (cpu_data_master_writedata),                                     //                                                     .writedata
		.cpu_data_master_debugaccess                                (cpu_data_master_debugaccess),                                   //                                                     .debugaccess
		.cpu_instruction_master_address                             (cpu_instruction_master_address),                                //                               cpu_instruction_master.address
		.cpu_instruction_master_waitrequest                         (cpu_instruction_master_waitrequest),                            //                                                     .waitrequest
		.cpu_instruction_master_read                                (cpu_instruction_master_read),                                   //                                                     .read
		.cpu_instruction_master_readdata                            (cpu_instruction_master_readdata),                               //                                                     .readdata
		.cpu_instruction_master_readdatavalid                       (cpu_instruction_master_readdatavalid),                          //                                                     .readdatavalid
		.audio_avalon_slave_address                                 (mm_interconnect_0_audio_avalon_slave_address),                  //                                   audio_avalon_slave.address
		.audio_avalon_slave_write                                   (mm_interconnect_0_audio_avalon_slave_write),                    //                                                     .write
		.audio_avalon_slave_read                                    (mm_interconnect_0_audio_avalon_slave_read),                     //                                                     .read
		.audio_avalon_slave_readdata                                (mm_interconnect_0_audio_avalon_slave_readdata),                 //                                                     .readdata
		.audio_avalon_slave_writedata                               (mm_interconnect_0_audio_avalon_slave_writedata),                //                                                     .writedata
		.cpu_jtag_debug_module_address                              (mm_interconnect_0_cpu_jtag_debug_module_address),               //                                cpu_jtag_debug_module.address
		.cpu_jtag_debug_module_write                                (mm_interconnect_0_cpu_jtag_debug_module_write),                 //                                                     .write
		.cpu_jtag_debug_module_read                                 (mm_interconnect_0_cpu_jtag_debug_module_read),                  //                                                     .read
		.cpu_jtag_debug_module_readdata                             (mm_interconnect_0_cpu_jtag_debug_module_readdata),              //                                                     .readdata
		.cpu_jtag_debug_module_writedata                            (mm_interconnect_0_cpu_jtag_debug_module_writedata),             //                                                     .writedata
		.cpu_jtag_debug_module_byteenable                           (mm_interconnect_0_cpu_jtag_debug_module_byteenable),            //                                                     .byteenable
		.cpu_jtag_debug_module_waitrequest                          (mm_interconnect_0_cpu_jtag_debug_module_waitrequest),           //                                                     .waitrequest
		.cpu_jtag_debug_module_debugaccess                          (mm_interconnect_0_cpu_jtag_debug_module_debugaccess),           //                                                     .debugaccess
		.cpu_peripheral_bridge_s0_address                           (mm_interconnect_0_cpu_peripheral_bridge_s0_address),            //                             cpu_peripheral_bridge_s0.address
		.cpu_peripheral_bridge_s0_write                             (mm_interconnect_0_cpu_peripheral_bridge_s0_write),              //                                                     .write
		.cpu_peripheral_bridge_s0_read                              (mm_interconnect_0_cpu_peripheral_bridge_s0_read),               //                                                     .read
		.cpu_peripheral_bridge_s0_readdata                          (mm_interconnect_0_cpu_peripheral_bridge_s0_readdata),           //                                                     .readdata
		.cpu_peripheral_bridge_s0_writedata                         (mm_interconnect_0_cpu_peripheral_bridge_s0_writedata),          //                                                     .writedata
		.cpu_peripheral_bridge_s0_burstcount                        (mm_interconnect_0_cpu_peripheral_bridge_s0_burstcount),         //                                                     .burstcount
		.cpu_peripheral_bridge_s0_byteenable                        (mm_interconnect_0_cpu_peripheral_bridge_s0_byteenable),         //                                                     .byteenable
		.cpu_peripheral_bridge_s0_readdatavalid                     (mm_interconnect_0_cpu_peripheral_bridge_s0_readdatavalid),      //                                                     .readdatavalid
		.cpu_peripheral_bridge_s0_waitrequest                       (mm_interconnect_0_cpu_peripheral_bridge_s0_waitrequest),        //                                                     .waitrequest
		.cpu_peripheral_bridge_s0_debugaccess                       (mm_interconnect_0_cpu_peripheral_bridge_s0_debugaccess),        //                                                     .debugaccess
		.DDR3_avl_address                                           (mm_interconnect_0_ddr3_avl_address),                            //                                             DDR3_avl.address
		.DDR3_avl_write                                             (mm_interconnect_0_ddr3_avl_write),                              //                                                     .write
		.DDR3_avl_read                                              (mm_interconnect_0_ddr3_avl_read),                               //                                                     .read
		.DDR3_avl_readdata                                          (mm_interconnect_0_ddr3_avl_readdata),                           //                                                     .readdata
		.DDR3_avl_writedata                                         (mm_interconnect_0_ddr3_avl_writedata),                          //                                                     .writedata
		.DDR3_avl_beginbursttransfer                                (mm_interconnect_0_ddr3_avl_beginbursttransfer),                 //                                                     .beginbursttransfer
		.DDR3_avl_burstcount                                        (mm_interconnect_0_ddr3_avl_burstcount),                         //                                                     .burstcount
		.DDR3_avl_byteenable                                        (mm_interconnect_0_ddr3_avl_byteenable),                         //                                                     .byteenable
		.DDR3_avl_readdatavalid                                     (mm_interconnect_0_ddr3_avl_readdatavalid),                      //                                                     .readdatavalid
		.DDR3_avl_waitrequest                                       (~mm_interconnect_0_ddr3_avl_waitrequest),                       //                                                     .waitrequest
		.jtag_uart_avalon_jtag_slave_address                        (mm_interconnect_0_jtag_uart_avalon_jtag_slave_address),         //                          jtag_uart_avalon_jtag_slave.address
		.jtag_uart_avalon_jtag_slave_write                          (mm_interconnect_0_jtag_uart_avalon_jtag_slave_write),           //                                                     .write
		.jtag_uart_avalon_jtag_slave_read                           (mm_interconnect_0_jtag_uart_avalon_jtag_slave_read),            //                                                     .read
		.jtag_uart_avalon_jtag_slave_readdata                       (mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata),        //                                                     .readdata
		.jtag_uart_avalon_jtag_slave_writedata                      (mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata),       //                                                     .writedata
		.jtag_uart_avalon_jtag_slave_waitrequest                    (mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest),     //                                                     .waitrequest
		.jtag_uart_avalon_jtag_slave_chipselect                     (mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect),      //                                                     .chipselect
		.onchip_memory2_1_s1_address                                (mm_interconnect_0_onchip_memory2_1_s1_address),                 //                                  onchip_memory2_1_s1.address
		.onchip_memory2_1_s1_write                                  (mm_interconnect_0_onchip_memory2_1_s1_write),                   //                                                     .write
		.onchip_memory2_1_s1_readdata                               (mm_interconnect_0_onchip_memory2_1_s1_readdata),                //                                                     .readdata
		.onchip_memory2_1_s1_writedata                              (mm_interconnect_0_onchip_memory2_1_s1_writedata),               //                                                     .writedata
		.onchip_memory2_1_s1_byteenable                             (mm_interconnect_0_onchip_memory2_1_s1_byteenable),              //                                                     .byteenable
		.onchip_memory2_1_s1_chipselect                             (mm_interconnect_0_onchip_memory2_1_s1_chipselect),              //                                                     .chipselect
		.onchip_memory2_1_s1_clken                                  (mm_interconnect_0_onchip_memory2_1_s1_clken),                   //                                                     .clken
		.spi_temperature_spi_control_port_address                   (mm_interconnect_0_spi_temperature_spi_control_port_address),    //                     spi_temperature_spi_control_port.address
		.spi_temperature_spi_control_port_write                     (mm_interconnect_0_spi_temperature_spi_control_port_write),      //                                                     .write
		.spi_temperature_spi_control_port_read                      (mm_interconnect_0_spi_temperature_spi_control_port_read),       //                                                     .read
		.spi_temperature_spi_control_port_readdata                  (mm_interconnect_0_spi_temperature_spi_control_port_readdata),   //                                                     .readdata
		.spi_temperature_spi_control_port_writedata                 (mm_interconnect_0_spi_temperature_spi_control_port_writedata),  //                                                     .writedata
		.spi_temperature_spi_control_port_chipselect                (mm_interconnect_0_spi_temperature_spi_control_port_chipselect), //                                                     .chipselect
		.sysid_qsys_control_slave_address                           (mm_interconnect_0_sysid_qsys_control_slave_address),            //                             sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata                          (mm_interconnect_0_sysid_qsys_control_slave_readdata),           //                                                     .readdata
		.timer_s1_address                                           (mm_interconnect_0_timer_s1_address),                            //                                             timer_s1.address
		.timer_s1_write                                             (mm_interconnect_0_timer_s1_write),                              //                                                     .write
		.timer_s1_readdata                                          (mm_interconnect_0_timer_s1_readdata),                           //                                                     .readdata
		.timer_s1_writedata                                         (mm_interconnect_0_timer_s1_writedata),                          //                                                     .writedata
		.timer_s1_chipselect                                        (mm_interconnect_0_timer_s1_chipselect)                          //                                                     .chipselect
	);

	audio_nios_mm_interconnect_1 mm_interconnect_1 (
		.altpll_outclk1_clk                                         (c2_out_clk_clk),                          //                                       altpll_outclk1.clk
		.cpu_peripheral_bridge_m0_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),          // cpu_peripheral_bridge_m0_reset_reset_bridge_in_reset.reset
		.key_reset_reset_bridge_in_reset_reset                      (rst_controller_003_reset_out_reset),      //                      key_reset_reset_bridge_in_reset.reset
		.cpu_peripheral_bridge_m0_address                           (cpu_peripheral_bridge_m0_address),        //                             cpu_peripheral_bridge_m0.address
		.cpu_peripheral_bridge_m0_waitrequest                       (cpu_peripheral_bridge_m0_waitrequest),    //                                                     .waitrequest
		.cpu_peripheral_bridge_m0_burstcount                        (cpu_peripheral_bridge_m0_burstcount),     //                                                     .burstcount
		.cpu_peripheral_bridge_m0_byteenable                        (cpu_peripheral_bridge_m0_byteenable),     //                                                     .byteenable
		.cpu_peripheral_bridge_m0_read                              (cpu_peripheral_bridge_m0_read),           //                                                     .read
		.cpu_peripheral_bridge_m0_readdata                          (cpu_peripheral_bridge_m0_readdata),       //                                                     .readdata
		.cpu_peripheral_bridge_m0_readdatavalid                     (cpu_peripheral_bridge_m0_readdatavalid),  //                                                     .readdatavalid
		.cpu_peripheral_bridge_m0_write                             (cpu_peripheral_bridge_m0_write),          //                                                     .write
		.cpu_peripheral_bridge_m0_writedata                         (cpu_peripheral_bridge_m0_writedata),      //                                                     .writedata
		.cpu_peripheral_bridge_m0_debugaccess                       (cpu_peripheral_bridge_m0_debugaccess),    //                                                     .debugaccess
		.i2c_scl_s1_address                                         (mm_interconnect_1_i2c_scl_s1_address),    //                                           i2c_scl_s1.address
		.i2c_scl_s1_write                                           (mm_interconnect_1_i2c_scl_s1_write),      //                                                     .write
		.i2c_scl_s1_readdata                                        (mm_interconnect_1_i2c_scl_s1_readdata),   //                                                     .readdata
		.i2c_scl_s1_writedata                                       (mm_interconnect_1_i2c_scl_s1_writedata),  //                                                     .writedata
		.i2c_scl_s1_chipselect                                      (mm_interconnect_1_i2c_scl_s1_chipselect), //                                                     .chipselect
		.i2c_sda_s1_address                                         (mm_interconnect_1_i2c_sda_s1_address),    //                                           i2c_sda_s1.address
		.i2c_sda_s1_write                                           (mm_interconnect_1_i2c_sda_s1_write),      //                                                     .write
		.i2c_sda_s1_readdata                                        (mm_interconnect_1_i2c_sda_s1_readdata),   //                                                     .readdata
		.i2c_sda_s1_writedata                                       (mm_interconnect_1_i2c_sda_s1_writedata),  //                                                     .writedata
		.i2c_sda_s1_chipselect                                      (mm_interconnect_1_i2c_sda_s1_chipselect), //                                                     .chipselect
		.key_s1_address                                             (mm_interconnect_1_key_s1_address),        //                                               key_s1.address
		.key_s1_write                                               (mm_interconnect_1_key_s1_write),          //                                                     .write
		.key_s1_readdata                                            (mm_interconnect_1_key_s1_readdata),       //                                                     .readdata
		.key_s1_writedata                                           (mm_interconnect_1_key_s1_writedata),      //                                                     .writedata
		.key_s1_chipselect                                          (mm_interconnect_1_key_s1_chipselect),     //                                                     .chipselect
		.pio_led_s1_address                                         (mm_interconnect_1_pio_led_s1_address),    //                                           pio_led_s1.address
		.pio_led_s1_write                                           (mm_interconnect_1_pio_led_s1_write),      //                                                     .write
		.pio_led_s1_readdata                                        (mm_interconnect_1_pio_led_s1_readdata),   //                                                     .readdata
		.pio_led_s1_writedata                                       (mm_interconnect_1_pio_led_s1_writedata),  //                                                     .writedata
		.pio_led_s1_chipselect                                      (mm_interconnect_1_pio_led_s1_chipselect), //                                                     .chipselect
		.sw_s1_address                                              (mm_interconnect_1_sw_s1_address),         //                                                sw_s1.address
		.sw_s1_write                                                (mm_interconnect_1_sw_s1_write),           //                                                     .write
		.sw_s1_readdata                                             (mm_interconnect_1_sw_s1_readdata),        //                                                     .readdata
		.sw_s1_writedata                                            (mm_interconnect_1_sw_s1_writedata),       //                                                     .writedata
		.sw_s1_chipselect                                           (mm_interconnect_1_sw_s1_chipselect)       //                                                     .chipselect
	);

	audio_nios_irq_mapper irq_mapper (
		.clk           (c0_001_out_clk_clk),                 //       clk.clk
		.reset         (rst_controller_002_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),           // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),           // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq),           // receiver2.irq
		.receiver3_irq (irq_mapper_receiver3_irq),           // receiver3.irq
		.receiver4_irq (irq_mapper_receiver4_irq),           // receiver4.irq
		.sender_irq    (cpu_d_irq_irq)                       //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer (
		.receiver_clk   (c2_out_clk_clk),                     //       receiver_clk.clk
		.sender_clk     (c0_001_out_clk_clk),                 //         sender_clk.clk
		.receiver_reset (rst_controller_003_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_002_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),      //           receiver.irq
		.sender_irq     (irq_mapper_receiver1_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_001 (
		.receiver_clk   (c2_out_clk_clk),                     //       receiver_clk.clk
		.sender_clk     (c0_001_out_clk_clk),                 //         sender_clk.clk
		.receiver_reset (rst_controller_003_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_002_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_001_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver2_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_002 (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (c0_001_out_clk_clk),                 //         sender_clk.clk
		.receiver_reset (rst_controller_008_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_002_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_002_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver3_irq)            //             sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (1)
	) irq_synchronizer_003 (
		.receiver_clk   (clk_clk),                            //       receiver_clk.clk
		.sender_clk     (c0_001_out_clk_clk),                 //         sender_clk.clk
		.receiver_reset (rst_controller_008_reset_out_reset), // receiver_clk_reset.reset
		.sender_reset   (rst_controller_002_reset_out_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_003_receiver_irq),  //           receiver.irq
		.sender_irq     (irq_mapper_receiver4_irq)            //             sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                 // reset_in0.reset
		.clk            (c2_out_clk_clk),                 //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_001 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (c0_001_out_clk_clk),                 //       clk.clk
		.reset_out      (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_002 (
		.reset_in0      (cpu_jtag_debug_module_reset_reset),      // reset_in0.reset
		.reset_in1      (~reset_reset_n),                         // reset_in1.reset
		.clk            (c0_001_out_clk_clk),                     //       clk.clk
		.reset_out      (rst_controller_002_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_002_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                                   // (terminated)
		.reset_req_in1  (1'b0),                                   // (terminated)
		.reset_in2      (1'b0),                                   // (terminated)
		.reset_req_in2  (1'b0),                                   // (terminated)
		.reset_in3      (1'b0),                                   // (terminated)
		.reset_req_in3  (1'b0),                                   // (terminated)
		.reset_in4      (1'b0),                                   // (terminated)
		.reset_req_in4  (1'b0),                                   // (terminated)
		.reset_in5      (1'b0),                                   // (terminated)
		.reset_req_in5  (1'b0),                                   // (terminated)
		.reset_in6      (1'b0),                                   // (terminated)
		.reset_req_in6  (1'b0),                                   // (terminated)
		.reset_in7      (1'b0),                                   // (terminated)
		.reset_req_in7  (1'b0),                                   // (terminated)
		.reset_in8      (1'b0),                                   // (terminated)
		.reset_req_in8  (1'b0),                                   // (terminated)
		.reset_in9      (1'b0),                                   // (terminated)
		.reset_req_in9  (1'b0),                                   // (terminated)
		.reset_in10     (1'b0),                                   // (terminated)
		.reset_req_in10 (1'b0),                                   // (terminated)
		.reset_in11     (1'b0),                                   // (terminated)
		.reset_req_in11 (1'b0),                                   // (terminated)
		.reset_in12     (1'b0),                                   // (terminated)
		.reset_req_in12 (1'b0),                                   // (terminated)
		.reset_in13     (1'b0),                                   // (terminated)
		.reset_req_in13 (1'b0),                                   // (terminated)
		.reset_in14     (1'b0),                                   // (terminated)
		.reset_req_in14 (1'b0),                                   // (terminated)
		.reset_in15     (1'b0),                                   // (terminated)
		.reset_req_in15 (1'b0)                                    // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_003 (
		.reset_in0      (cpu_jtag_debug_module_reset_reset),  // reset_in0.reset
		.reset_in1      (~reset_reset_n),                     // reset_in1.reset
		.clk            (c2_out_clk_clk),                     //       clk.clk
		.reset_out      (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_004 (
		.reset_in0      (cpu_jtag_debug_module_reset_reset),  // reset_in0.reset
		.reset_in1      (~reset_reset_n),                     // reset_in1.reset
		.clk            (c0_out_clk_clk),                     //       clk.clk
		.reset_out      (rst_controller_004_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_005 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_005_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_006 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_006_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("none"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_007 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.clk            (),                                   //       clk.clk
		.reset_out      (rst_controller_007_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_008 (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (cpu_jtag_debug_module_reset_reset),  // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_008_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller_009 (
		.reset_in0      (~ddr3_afi_reset_reset),              // reset_in0.reset
		.clk            (ddr3_afi_clk_clk),                   //       clk.clk
		.reset_out      (rst_controller_009_reset_out_reset), // reset_out.reset
		.reset_req      (),                                   // (terminated)
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_in1      (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
